module wallace_tree_24x24 (
    input  [23:0] a,
    input  [23:0] b,
    output [47:8] x,  //sum high
    output [47:8] y,  //carry high
    output [ 7:0] z   //sum low

);
  parameter zero = 1'b0;
  reg [23:00] a_b [23:00];
  integer i, j;

  always @(*) begin
    for (i = 0; i < 24; i = i + 1)
      for (j = 0; j < 24; j = j + 1)
        a_b[i][j] = a[i] & b[j];
  end

  //--------------------------------------------------------------------------------
 
  wire [7:0] s1 [44:1];
  wire [7:0] c1 [45:2];

  full_adder l1_01_1(a_b[00][01],a_b[01][00],zero,s1[01][00],c1[02][00]); // l1 means layer 1 , s[01] 01 means the bit seq num , 1 means the seq of full_adder 
                                                                         // c1[02] 02 means the bit seq num of full_adder that c1 will connect
  full_adder l1_02_1(a_b[00][02],a_b[01][01],a_b[02][00],s1[02][00],c1[03][00]);

  full_adder l1_03_1(a_b[00][03],a_b[01][02],a_b[02][01],s1[03][00],c1[04][00]);// [03][00] connect to layer2

  full_adder l1_04_1(a_b[00][04],a_b[01][03],a_b[02][02],s1[04][00],c1[05][00]);
  full_adder l1_04_2(a_b[03][01],a_b[04][00],zero,s1[04][01],c1[05][01]); 
  //c1[05][01] to layer3
  //layer2 与 layer1 直接同列的csa存在数量差，进位插到下层去，同位不用担心，有
  //三个输入位能处理同位的数据

  full_adder l1_05_1(a_b[00][05],a_b[01][04],a_b[02][03],s1[05][00],c1[06][00]);
  full_adder l1_05_2(a_b[03][02],a_b[04][01],a_b[05][00],s1[05][01],c1[06][01]);

  full_adder l1_06_1(a_b[00][06],a_b[01][05],a_b[02][04],s1[06][00],c1[07][00]);
  full_adder l1_06_2(a_b[03][03],a_b[04][02],a_b[05][01],s1[06][01],c1[07][01]); // [06][00] connect to layer2

  genvar k;

  generate
    for (k = 0 ; k < 2; k = k+1) begin: l1_07
      full_adder l1_07(a_b[3*k][07-3*k],a_b[3*k+1][7-3*k-1],a_b[3*k+2][7-3*k-2],s1[07][k],c1[08][k]);
    end
  endgenerate

      full_adder l1_07_2(a_b[06][01],a_b[07][00],zero,s1[07][02],c1[08][02]);

  generate
    for (k = 0 ; k < 3; k = k+1) begin: l1_08
      full_adder l1_08(a_b[3*k][08-3*k],a_b[3*k+1][8-3*k-1],a_b[3*k+2][8-3*k-2],s1[08][k],c1[09][k]);
    end
  endgenerate

  generate
    for (k = 0 ; k < 3; k = k+1) begin: l1_09
      full_adder l1_09(a_b[3*k][09-3*k],a_b[3*k+1][9-3*k-1],a_b[3*k+2][9-3*k-2],s1[09][k],c1[10][k]);
    end
  endgenerate // [09][00] connect to layer2

  generate
    for (k = 0 ; k < 3; k = k+1) begin: l1_10
      full_adder l1_10(a_b[3*k][10-3*k],a_b[3*k+1][10-3*k-1],a_b[3*k+2][10-3*k-2],s1[10][k],c1[11][k]);
    end
  endgenerate

      full_adder l1_10_3(a_b[09][01],a_b[10][00],zero,s1[10][03],c1[11][03]);

  generate
    for (k = 0 ; k < 4; k = k+1) begin: l1_11
      full_adder l1_11(a_b[3*k][11-3*k],a_b[3*k+1][11-3*k-1],a_b[3*k+2][11-3*k-2],s1[11][k],c1[12][k]);
    end
  endgenerate

  generate
    for (k = 0 ; k < 4; k = k+1) begin: l1_12
      full_adder l1_12(a_b[3*k][12-3*k],a_b[3*k+1][12-3*k-1],a_b[3*k+2][12-3*k-2],s1[12][k],c1[13][k]);
    end
  endgenerate // [12][00] connect to layer2

  generate
    for (k = 0 ; k < 4; k = k+1) begin: l1_13
      full_adder l1_13(a_b[3*k][13-3*k],a_b[3*k+1][13-3*k-1],a_b[3*k+2][13-3*k-2],s1[13][k],c1[14][k]);
    end
  endgenerate

      full_adder l1_13_4(a_b[12][01],a_b[13][00],zero,s1[13][4],c1[14][4]);

  generate
    for (k = 0 ; k < 5; k = k+1) begin: l1_14
      full_adder l1_14(a_b[3*k][14-3*k],a_b[3*k+1][14-3*k-1],a_b[3*k+2][14-3*k-2],s1[14][k],c1[15][k]);
    end
  endgenerate

  generate
    for (k = 0 ; k < 5; k = k+1) begin: l1_15
      full_adder l1_15(a_b[3*k][15-3*k],a_b[3*k+1][15-3*k-1],a_b[3*k+2][15-3*k-2],s1[15][k],c1[16][k]);
    end
  endgenerate // [15][00]

  generate
    for (k = 0 ; k < 5; k = k+1) begin: l1_16
      full_adder l1_16(a_b[3*k][16-3*k],a_b[3*k+1][16-3*k-1],a_b[3*k+2][16-3*k-2],s1[16][k],c1[17][k]);
    end
  endgenerate

      full_adder l1_16_5(a_b[15][1],a_b[16][0],zero,s1[16][5],c1[17][5]);

  generate
    for (k = 0 ; k < 6; k = k+1) begin: l1_17
      full_adder l1_17(a_b[3*k][17-3*k],a_b[3*k+1][17-3*k-1],a_b[3*k+2][17-3*k-2],s1[17][k],c1[18][k]);
    end
  endgenerate

  generate
    for (k = 0 ; k < 6; k = k+1) begin: l1_18
      full_adder l1_18(a_b[3*k][18-3*k],a_b[3*k+1][18-3*k-1],a_b[3*k+2][18-3*k-2],s1[18][k],c1[19][k]);
    end
  endgenerate // [18][00] connect to layer2

  generate
    for (k = 0 ; k < 6; k = k+1) begin: l1_19
      full_adder l1_19(a_b[3*k][19-3*k],a_b[3*k+1][19-3*k-1],a_b[3*k+2][19-3*k-2],s1[19][k],c1[20][k]);
    end
  endgenerate 
      full_adder l1_19_6(a_b[18][1],a_b[19][0],zero,s1[19][6],c1[20][6]);

  generate
    for (k = 0 ; k < 7; k = k+1) begin: l1_20
      full_adder l1_20(a_b[3*k][20-3*k],a_b[3*k+1][20-3*k-1],a_b[3*k+2][20-3*k-2],s1[20][k],c1[21][k]);
    end
  endgenerate 

  generate
    for (k = 0 ; k < 7; k = k+1) begin: l1_21
      full_adder l1_21(a_b[3*k][21-3*k],a_b[3*k+1][21-3*k-1],a_b[3*k+2][21-3*k-2],s1[21][k],c1[22][k]);
    end
  endgenerate // [21][00] connect to layer2

  generate
    for (k = 0 ; k < 7; k = k+1) begin: l1_22
      full_adder l1_22(a_b[3*k][22-3*k],a_b[3*k+1][22-3*k-1],a_b[3*k+2][22-3*k-2],s1[22][k],c1[23][k]);
    end
  endgenerate

      full_adder l1_22_7(a_b[21][1],a_b[22][0],zero,s1[22][7],c1[23][7]);

  generate
    for (k = 0 ; k < 8; k = k+1) begin: l1_23
      full_adder l1_23(a_b[3*k][23-3*k],a_b[3*k+1][23-3*k-1],a_b[3*k+2][23-3*k-2],s1[23][k],c1[24][k]);
    end
  endgenerate

  generate
    for (k = 0 ; k < 7; k = k+1) begin: l1_24
      full_adder l1_24(a_b[23-3*k][3*k+1],a_b[23-3*k-1][3*k+2],a_b[23-3*k-2][3*k+3],s1[24][k],c1[25][k]);
    end
  endgenerate

      full_adder l1_24_7(a_b[02][22],a_b[01][23],zero,s1[24][7],c1[25][7]);

  generate
    for (k = 0 ; k < 7; k = k+1) begin: l1_25
      full_adder l1_25(a_b[23-3*k][3*k+2],a_b[23-3*k-1][3*k+3],a_b[23-3*k-2][3*k+4],s1[25][k],c1[26][k]);
    end
  endgenerate // [2][23] connect to layer2

  generate
    for (k = 0 ; k < 7; k = k+1) begin: l1_26
      full_adder l1_26(a_b[23-3*k][3*k+3],a_b[23-3*k-1][3*k+4],a_b[23-3*k-2][3*k+5],s1[26][k],c1[27][k]);
    end
  endgenerate

  generate
    for (k = 0 ; k < 6; k = k+1) begin: l1_27
      full_adder l1_27(a_b[23-3*k][3*k+4],a_b[23-3*k-1][3*k+5],a_b[23-3*k-2][3*k+6],s1[27][k],c1[28][k]);
    end
  endgenerate

      full_adder l1_27_6(a_b[05][22],a_b[04][23],zero,s1[27][6],c1[28][6]);

  generate
    for (k = 0 ; k < 6; k = k+1) begin: l1_28
      full_adder l1_28(a_b[23-3*k][3*k+5],a_b[23-3*k-1][3*k+6],a_b[23-3*k-2][3*k+7],s1[28][k],c1[29][k]);
    end
  endgenerate //[5][23] connect to layer2

  generate
    for (k = 0 ; k < 6; k = k+1) begin: l1_29
      full_adder l1_29(a_b[23-3*k][3*k+6],a_b[23-3*k-1][3*k+7],a_b[23-3*k-2][3*k+8],s1[29][k],c1[30][k]);
    end
  endgenerate 

  generate
    for (k = 0 ; k < 5; k = k+1) begin: l1_30
      full_adder l1_30(a_b[23-3*k][3*k+7],a_b[23-3*k-1][3*k+8],a_b[23-3*k-2][3*k+9],s1[30][k],c1[31][k]);
    end
  endgenerate 

      full_adder l1_30_5(a_b[08][22],a_b[07][23],zero,s1[30][5],c1[31][5]);

  generate
    for (k = 0 ; k < 5; k = k+1) begin: l1_31
      full_adder l1_31(a_b[23-3*k][3*k+8],a_b[23-3*k-1][3*k+9],a_b[23-3*k-2][3*k+10],s1[31][k],c1[32][k]);
    end
  endgenerate // [8][23] connect to layer2

  generate
    for (k = 0 ; k < 5; k = k+1) begin: l1_32
      full_adder l1_32(a_b[23-3*k][3*k+9],a_b[23-3*k-1][3*k+10],a_b[23-3*k-2][3*k+11],s1[32][k],c1[33][k]);
    end
  endgenerate 

  generate
    for (k = 0 ; k < 4; k = k+1) begin: l1_33
      full_adder l1_33(a_b[23-3*k][3*k+10],a_b[23-3*k-1][3*k+11],a_b[23-3*k-2][3*k+12],s1[33][k],c1[34][k]);
    end
  endgenerate 

      full_adder l1_33_4(a_b[11][22],a_b[10][23],zero,s1[33][4],c1[34][4]);

  generate
    for (k = 0 ; k < 4; k = k+1) begin: l1_34
      full_adder l1_34(a_b[23-3*k][3*k+11],a_b[23-3*k-1][3*k+12],a_b[23-3*k-2][3*k+13],s1[34][k],c1[35][k]);
    end
  endgenerate //[11][23] connect to layer2

  generate
    for (k = 0 ; k < 4; k = k+1) begin: l1_35
      full_adder l1_35(a_b[23-3*k][3*k+12],a_b[23-3*k-1][3*k+13],a_b[23-3*k-2][3*k+14],s1[35][k],c1[36][k]);
    end
  endgenerate

  generate
    for (k = 0 ; k < 3; k = k+1) begin: l1_36
      full_adder l1_36(a_b[23-3*k][3*k+13],a_b[23-3*k-1][3*k+14],a_b[23-3*k-2][3*k+15],s1[36][k],c1[37][k]);
    end
  endgenerate

      full_adder l1_36_3(a_b[14][22],a_b[13][23],zero,s1[36][3],c1[37][3]);

      full_adder l1_44(a_b[21][23],a_b[22][22],a_b[23][21],s1[44][0],c1[45][0]);

      full_adder l1_43(a_b[21][22],a_b[22][21],a_b[23][20],s1[43][0],c1[44][0]);// [20][23] connect to layer2

      full_adder l1_42_1(a_b[21][21],a_b[22][20],a_b[23][19],s1[42][0],c1[43][0]);
      full_adder l1_42_2(a_b[20][22],a_b[19][23],zero,s1[42][1],c1[43][1]);

      full_adder l1_41_1(a_b[21][20],a_b[22][19],a_b[23][18],s1[41][0],c1[42][0]);
      full_adder l1_41_2(a_b[20][21],a_b[19][22],a_b[18][23],s1[41][1],c1[42][1]);

      full_adder l1_40_1(a_b[21][19],a_b[22][18],a_b[23][17],s1[40][0],c1[41][0]);
      full_adder l1_40_2(a_b[20][20],a_b[19][21],a_b[18][22],s1[40][1],c1[41][1]);// [17][23] connect to layer2

      full_adder l1_39_1(a_b[21][18],a_b[22][17],a_b[23][16],s1[39][0],c1[40][0]);
      full_adder l1_39_2(a_b[20][19],a_b[19][20],a_b[18][21],s1[39][1],c1[40][1]);
      full_adder l1_39_3(a_b[17][22],a_b[16][23],zero,s1[39][2],c1[40][2]);

      full_adder l1_38_1(a_b[21][17],a_b[22][16],a_b[23][15],s1[38][0],c1[39][0]);
      full_adder l1_38_2(a_b[20][18],a_b[19][19],a_b[18][20],s1[38][1],c1[39][1]);
      full_adder l1_38_3(a_b[17][21],a_b[16][22],a_b[15][23],s1[38][2],c1[39][2]);

      full_adder l1_37_1(a_b[21][16],a_b[22][15],a_b[23][14],s1[37][0],c1[38][0]);
      full_adder l1_37_2(a_b[20][17],a_b[19][18],a_b[18][19],s1[37][1],c1[38][1]);
      full_adder l1_37_3(a_b[17][20],a_b[16][21],a_b[15][22],s1[37][2],c1[38][2]);// [14][23] connect to layer2


  //level1--------------------------------------------------------------------------


  //level2--------------------------------------------------------------------------
 
  wire [4:0] s2[45:2];
  wire [4:0] c2[46:3];

  full_adder l2_02(s1[02][00],c1[02][00],zero,s2[02][00],c2[03][00]);

  full_adder l2_03(s1[03][00],c1[03][00],a_b[03][00],s2[03][00],c2[04][00]);

  full_adder l2_04(s1[04][00],c1[04][00],s1[04][01],s2[04][00],c2[05][00]);

  full_adder l2_05(s1[05][00],c1[05][00],s1[05][01],s2[05][00],c2[06][00]);
  //c1[05][01] to layer3

  full_adder l2_06_1(s1[06][00],c1[06][00],a_b[06][00],s2[06][00],c2[07][00]);
  full_adder l2_06_2(s1[06][01],c1[06][01],zero,s2[06][01],c2[07][01]);

  full_adder l2_07_1(s1[07][00],c1[07][00],zero,s2[07][00],c2[08][00]);
  full_adder l2_07_2(s1[07][01],c1[07][01],s1[07][02],s2[07][01],c2[08][01]);

  full_adder l2_08_1(s1[08][00],c1[08][00],c1[08][02],s2[08][00],c2[09][00]);
  full_adder l2_08_2(s1[08][01],c1[08][01],s1[08][02],s2[08][01],c2[09][01]);

  full_adder l2_09_1(s1[09][00],s1[09][01],s1[09][02],s2[09][00],c2[10][00]);
  full_adder l2_09_2(a_b[09][00],c1[09][01],c1[09][02],s2[09][01],c2[10][01]);
  //c1[09][00] to layer3

  full_adder l2_10_1(s1[10][00],s1[10][01],s1[10][02],s2[10][00],c2[11][00]);
  full_adder l2_10_2(s1[10][03],c1[10][01],c1[10][02],s2[10][01],c2[11][01]);
  //c1[10][00] to layer3

  full_adder l2_11_1(s1[11][00],s1[11][01],s1[11][02],s2[11][00],c2[12][00]);
  full_adder l2_11_2(s1[11][03],c1[11][00],c1[11][01],s2[11][01],c2[12][01]);
  full_adder l2_11_3(c1[11][02],c1[11][03],zero,s2[11][02],c2[12][02]);

  full_adder l2_12_1(s1[12][00],s1[12][01],s1[12][02],s2[12][00],c2[13][00]);
  full_adder l2_12_2(s1[12][03],c1[12][00],c1[12][01],s2[12][01],c2[13][01]);
  full_adder l2_12_3(c1[12][02],c1[12][03],a_b[12][00],s2[12][02],c2[13][02]);

  full_adder l2_13_1(s1[13][00],s1[13][01],s1[13][02],s2[13][00],c2[14][00]);
  full_adder l2_13_2(s1[13][03],s1[13][04],c1[13][00],s2[13][01],c2[14][01]);
  full_adder l2_13_3(c1[13][01],c1[13][02],c1[13][03],s2[13][02],c2[14][02]);

  full_adder l2_14_1(s1[14][00],s1[14][01],s1[14][02],s2[14][00],c2[15][00]);
  full_adder l2_14_2(s1[14][03],s1[14][04],c1[14][04],s2[14][01],c2[15][01]);
  full_adder l2_14_3(c1[14][01],c1[14][02],c1[14][03],s2[14][02],c2[15][02]);
  //c1[14][00] to layer3
  
  full_adder l2_15_1(s1[15][00],s1[15][01],s1[15][02],s2[15][00],c2[16][00]);
  full_adder l2_15_2(s1[15][03],s1[15][04],c1[15][00],s2[15][01],c2[16][01]);
  full_adder l2_15_3(c1[15][01],c1[15][02],c1[15][03],s2[15][02],c2[16][02]);
  full_adder l2_15_4(c1[15][04],a_b[15][00],zero,s2[15][03],c2[16][03]);

  full_adder l2_16_1(s1[16][00],s1[16][01],s1[16][02],s2[16][00],c2[17][00]);
  full_adder l2_16_2(s1[16][03],s1[16][04],s1[16][05],s2[16][01],c2[17][01]);
  full_adder l2_16_3(c1[16][00],c1[16][01],c1[16][02],s2[16][02],c2[17][02]);
  full_adder l2_16_4(c1[16][03],c1[16][04],zero,s2[16][03],c2[17][03]);

  full_adder l2_17_1(s1[17][00],s1[17][01],s1[17][02],s2[17][00],c2[18][00]);
  full_adder l2_17_2(s1[17][03],s1[17][04],s1[17][05],s2[17][01],c2[18][01]);
  full_adder l2_17_3(c1[17][00],c1[17][01],c1[17][02],s2[17][02],c2[18][02]);
  full_adder l2_17_4(c1[17][03],c1[17][04],c1[17][05],s2[17][03],c2[18][03]);

  full_adder l2_18_1(s1[18][00],s1[18][01],s1[18][02],s2[18][00],c2[19][00]);
  full_adder l2_18_2(s1[18][03],s1[18][04],s1[18][05],s2[18][01],c2[19][01]);
  full_adder l2_18_3(a_b[18][00],c1[18][01],c1[18][02],s2[18][02],c2[19][02]);
  full_adder l2_18_4(c1[18][03],c1[18][04],c1[18][05],s2[18][03],c2[19][03]);
  //c1[18][00] to layer3
  //

  full_adder l2_19_1(s1[19][00],s1[19][01],s1[19][02],s2[19][00],c2[20][00]);
  full_adder l2_19_2(s1[19][03],s1[19][04],s1[19][05],s2[19][01],c2[20][01]);
  full_adder l2_19_3(s1[19][06],c1[19][01],c1[19][02],s2[19][02],c2[20][02]);
  full_adder l2_19_4(c1[19][03],c1[19][04],c1[19][05],s2[19][03],c2[20][03]);
  //c1[19][00] to layer3
  //
  full_adder l2_20_1(s1[20][00],s1[20][01],s1[20][02],s2[20][00],c2[21][00]);
  full_adder l2_20_2(s1[20][03],s1[20][04],s1[20][05],s2[20][01],c2[21][01]);
  full_adder l2_20_3(s1[20][06],c1[20][01],c1[20][02],s2[20][02],c2[21][02]);
  full_adder l2_20_4(c1[20][03],c1[20][04],c1[20][05],s2[20][03],c2[21][03]);
  full_adder l2_20_5(c1[20][06],c1[20][00],zero,s2[20][04],c2[21][04]);

  full_adder l2_21_1(s1[21][00],s1[21][01],s1[21][02],s2[21][00],c2[22][00]);
  full_adder l2_21_2(s1[21][03],s1[21][04],s1[21][05],s2[21][01],c2[22][01]);
  full_adder l2_21_3(s1[21][06],c1[21][01],c1[21][02],s2[21][02],c2[22][02]);
  full_adder l2_21_4(c1[21][03],c1[21][04],c1[21][05],s2[21][03],c2[22][03]);
  full_adder l2_21_5(c1[21][06],c1[21][00],a_b[21][00],s2[21][04],c2[22][04]);

  full_adder l2_22_1(s1[22][00],s1[22][01],s1[22][02],s2[22][00],c2[23][00]);
  full_adder l2_22_2(s1[22][03],s1[22][04],s1[22][05],s2[22][01],c2[23][01]);
  full_adder l2_22_3(s1[22][06],s1[22][07],c1[22][00],s2[22][02],c2[23][02]);
  full_adder l2_22_4(c1[22][01],c1[22][02],c1[22][03],s2[22][03],c2[23][03]);
  full_adder l2_22_5(c1[22][04],c1[22][05],c1[22][06],s2[22][04],c2[23][04]);

  full_adder l2_23_1(s1[23][00],s1[23][01],s1[23][02],s2[23][00],c2[24][00]);
  full_adder l2_23_2(s1[23][03],s1[23][04],s1[23][05],s2[23][01],c2[24][01]);
  full_adder l2_23_3(s1[23][06],s1[23][07],c1[23][00],s2[23][02],c2[24][02]);
  full_adder l2_23_4(c1[23][01],c1[23][02],c1[23][03],s2[23][03],c2[24][03]);
  full_adder l2_23_5(c1[23][04],c1[23][05],c1[23][06],s2[23][04],c2[24][04]);
  // c1[23][7] to layer3
  full_adder l2_24_1(s1[24][00],s1[24][01],s1[24][02],s2[24][00],c2[25][00]);
  full_adder l2_24_2(s1[24][03],s1[24][04],s1[24][05],s2[24][01],c2[25][01]);
  full_adder l2_24_3(s1[24][06],s1[24][07],c1[24][00],s2[24][02],c2[25][02]);
  full_adder l2_24_4(c1[24][01],c1[24][02],c1[24][03],s2[24][03],c2[25][03]);
  full_adder l2_24_5(c1[24][04],c1[24][05],c1[24][06],s2[24][04],c2[25][04]);
  // c1[24][7] to layer3
  full_adder l2_25_1(s1[25][00],s1[25][01],s1[25][02],s2[25][00],c2[26][00]);
  full_adder l2_25_2(s1[25][03],s1[25][04],s1[25][05],s2[25][01],c2[26][01]);
  full_adder l2_25_3(s1[25][06],a_b[2][23],c1[25][00],s2[25][02],c2[26][02]);
  full_adder l2_25_4(c1[25][01],c1[25][02],c1[25][03],s2[25][03],c2[26][03]);
  full_adder l2_25_5(c1[25][04],c1[25][05],c1[25][06],s2[25][04],c2[26][04]);
  // c1[25][7] to layer3
  
  full_adder l2_26_1(s1[26][00],s1[26][01],s1[26][02],s2[26][00],c2[27][00]);
  full_adder l2_26_2(s1[26][03],s1[26][04],s1[26][05],s2[26][01],c2[27][01]);
  full_adder l2_26_3(s1[26][06],zero,c1[26][00],s2[26][02],c2[27][02]);
  full_adder l2_26_4(c1[26][01],c1[26][02],c1[26][03],s2[26][03],c2[27][03]);
  full_adder l2_26_5(c1[26][04],c1[26][05],c1[26][06],s2[26][04],c2[27][04]);

  full_adder l2_27_1(s1[27][00],s1[27][01],s1[27][02],s2[27][00],c2[28][00]);
  full_adder l2_27_2(s1[27][03],s1[27][04],s1[27][05],s2[27][01],c2[28][01]);
  full_adder l2_27_3(s1[27][06],zero,c1[27][00],s2[27][02],c2[28][02]);
  full_adder l2_27_4(c1[27][01],c1[27][02],c1[27][03],s2[27][03],c2[28][03]);
  full_adder l2_27_5(c1[27][04],c1[27][05],c1[27][06],s2[27][04],c2[28][04]);

  full_adder l2_28_1(s1[28][00],s1[28][01],s1[28][02],s2[28][00],c2[29][00]);
  full_adder l2_28_2(s1[28][03],s1[28][04],s1[28][05],s2[28][01],c2[29][01]);
  full_adder l2_28_3(a_b[5][23],zero,c1[28][00],s2[28][02],c2[29][02]);
  full_adder l2_28_4(c1[28][01],c1[28][02],c1[28][03],s2[28][03],c2[29][03]);
  full_adder l2_28_5(c1[28][04],c1[28][05],c1[28][06],s2[28][04],c2[29][04]);

  full_adder l2_29_1(s1[29][00],s1[29][01],s1[29][02],s2[29][00],c2[30][00]);
  full_adder l2_29_2(s1[29][03],s1[29][04],s1[29][05],s2[29][01],c2[30][01]);
  full_adder l2_29_3(c1[29][00],c1[29][01],c1[29][02],s2[29][02],c2[30][02]);
  full_adder l2_29_4(c1[29][03],c1[29][04],c1[29][05],s2[29][03],c2[30][03]);

  full_adder l2_30_1(s1[30][00],s1[30][01],s1[30][02],s2[30][00],c2[31][00]);
  full_adder l2_30_2(s1[30][03],s1[30][04],s1[30][05],s2[30][01],c2[31][01]);
  full_adder l2_30_3(c1[30][00],c1[30][01],c1[30][02],s2[30][02],c2[31][02]);
  full_adder l2_30_4(c1[30][03],c1[30][04],c1[30][05],s2[30][03],c2[31][03]);

  full_adder l2_31_1(s1[31][00],s1[31][01],s1[31][02],s2[31][00],c2[32][00]);
  full_adder l2_31_2(s1[31][03],s1[31][04],a_b[8][23],s2[31][01],c2[32][01]);
  full_adder l2_31_3(c1[31][00],c1[31][01],c1[31][02],s2[31][02],c2[32][02]);
  full_adder l2_31_4(c1[31][03],c1[31][04],c1[31][05],s2[31][03],c2[32][03]);

  full_adder l2_32_1(s1[32][00],s1[32][01],s1[32][02],s2[32][00],c2[33][00]);
  full_adder l2_32_2(s1[32][03],s1[32][04],c1[32][03],s2[32][01],c2[33][01]);
  full_adder l2_32_3(c1[32][00],c1[32][01],c1[32][02],s2[32][02],c2[33][02]);
  // c1[32][04] to layer3
  full_adder l2_33_1(s1[33][00],s1[33][01],s1[33][02],s2[33][00],c2[34][00]);
  full_adder l2_33_2(s1[33][03],s1[33][04],c1[33][03],s2[33][01],c2[34][01]);
  full_adder l2_33_3(c1[33][00],c1[33][01],c1[33][02],s2[33][02],c2[34][02]);
  // c1[33][04] to layer3
  full_adder l2_34_1(s1[34][00],s1[34][01],s1[34][02],s2[34][00],c2[35][00]);
  full_adder l2_34_2(s1[34][03],a_b[11][23],c1[34][03],s2[34][01],c2[35][01]);
  full_adder l2_34_3(c1[34][00],c1[34][01],c1[34][02],s2[34][02],c2[35][02]);
  // c1[34][04] to layer3

  full_adder l2_35_1(s1[35][00],s1[35][01],s1[35][02],s2[35][00],c2[36][00]);
  full_adder l2_35_2(s1[35][03],zero,c1[35][03],s2[35][01],c2[36][01]);
  full_adder l2_35_3(c1[35][00],c1[35][01],c1[35][02],s2[35][02],c2[36][02]);

  full_adder l2_36_1(s1[36][00],s1[36][01],s1[36][02],s2[36][00],c2[37][00]);
  full_adder l2_36_2(s1[36][03],zero,c1[36][03],s2[36][01],c2[37][01]);
  full_adder l2_36_3(c1[36][00],c1[36][01],c1[36][02],s2[36][02],c2[37][02]);

  full_adder l2_37_1(s1[37][00],s1[37][01],s1[37][02],s2[37][00],c2[38][00]);
  full_adder l2_37_2(a_b[14][23],zero,c1[37][03],s2[37][01],c2[38][01]);
  full_adder l2_37_3(c1[37][00],c1[37][01],c1[37][02],s2[37][02],c2[38][02]);

  full_adder l2_38_1(s1[38][00],s1[38][01],s1[38][02],s2[38][00],c2[39][00]);
  full_adder l2_38_2(c1[38][00],c1[38][01],c1[38][02],s2[38][01],c2[39][01]);

  full_adder l2_39_1(s1[39][00],s1[39][01],s1[39][02],s2[39][00],c2[40][00]);
  full_adder l2_39_2(c1[39][00],c1[39][01],c1[39][02],s2[39][01],c2[40][01]);

  full_adder l2_40_1(s1[40][00],s1[40][01],a_b[17][23],s2[40][00],c2[41][00]);
  full_adder l2_40_2(c1[40][00],c1[40][01],c1[40][02],s2[40][01],c2[41][01]);

  full_adder l2_41_1(s1[41][00],s1[41][01],c1[41][00],s2[41][00],c2[42][00]);
  // c1[41][1] to layer3
  
  full_adder l2_42_1(s1[42][00],s1[42][01],c1[42][00],s2[42][00],c2[43][00]);
  // c1[42][1] to layer3
  
  full_adder l2_43_1(s1[43][00],a_b[20][23],c1[43][00],s2[43][00],c2[44][00]);
  // c1[43][1] to layer3

  full_adder l2_44_1(s1[44][00],zero,c1[44][00],s2[44][00],c2[45][00]);

  full_adder l2_45_1(a_b[23][22],a_b[22][23],c1[45][00],s2[45][00],c2[46][00]);
  //level2--------------------------------------------------------------------------
  
  wire [3:0] s3[43:3];
  wire [3:0] c3[44:4];

  full_adder l3_03_1(s2[03][00],c2[03][00],zero,s3[03][00],c3[04][00]);

  full_adder l3_04_1(s2[04][00],c2[04][00],zero,s3[04][00],c3[05][00]);

  full_adder l3_05_1(s2[05][00],c2[05][00],c1[05][01],s3[05][00],c3[06][00]);

  full_adder l3_06_1(s2[06][00],c2[06][00],zero,s3[06][00],c3[07][00]);

  full_adder l3_07_1(s2[07][00],s2[07][01],c2[07][00],s3[07][00],c3[08][00]);
  // c2[07][01] to layer4
  full_adder l3_08_1(s2[08][00],s2[08][01],c2[08][00],s3[08][00],c3[09][00]);
  // c2[08][01] to layer4
  
  //level3--------------------------------------------------------------------------

  assign z[0] = a_b[0][0];
  assign z[1] = s1[01][00];
  assign z[2] = s2[02][00];

endmodule

