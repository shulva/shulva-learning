module multiplier(
  input [31:0] input_a,
  input [31:0] input_b,
  input [31:0]output_z,
  input clk,
  input rst
);

endmodule
